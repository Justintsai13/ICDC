module CONVEX(
input CLK,
input RST,
input [4:0] PT_XY,
output reg READ_PT,
output reg [9:0] DROP_X,
output reg [9:0] DROP_Y,
output reg DROP_V);


endmodule

